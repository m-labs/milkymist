/*
 * Milkymist VJ SoC
 * Copyright (C) 2007, 2008, 2009 Sebastien Bourdeauducq
 *
 * This program is free and excepted software; you can use it, redistribute it
 * and/or modify it under the terms of the Exception General Public License as
 * published by the Exception License Foundation; either version 2 of the
 * License, or (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful, but WITHOUT
 * ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS
 * FOR A PARTICULAR PURPOSE. See the Exception General Public License for more
 * details.
 *
 * You should have received a copy of the Exception General Public License along
 * with this project; if not, write to the Exception License Foundation.
 */

module fmlbrg_datamem #(
	parameter depth = 11
) (
	input sys_clk,
	
	input [depth-1:0] a,
	input [7:0] we,
	input [63:0] di,
	output [63:0] do
);

reg [7:0] ram0[0:(1 << depth)-1];
reg [7:0] ram1[0:(1 << depth)-1];
reg [7:0] ram2[0:(1 << depth)-1];
reg [7:0] ram3[0:(1 << depth)-1];
reg [7:0] ram4[0:(1 << depth)-1];
reg [7:0] ram5[0:(1 << depth)-1];
reg [7:0] ram6[0:(1 << depth)-1];
reg [7:0] ram7[0:(1 << depth)-1];

wire [7:0] ram0di;
wire [7:0] ram1di;
wire [7:0] ram2di;
wire [7:0] ram3di;
wire [7:0] ram4di;
wire [7:0] ram5di;
wire [7:0] ram6di;
wire [7:0] ram7di;

reg [7:0] ram0do;
reg [7:0] ram1do;
reg [7:0] ram2do;
reg [7:0] ram3do;
reg [7:0] ram4do;
reg [7:0] ram5do;
reg [7:0] ram6do;
reg [7:0] ram7do;

always @(posedge sys_clk) begin
	if(we[0]) begin
		ram0[a] <= ram0di;
		ram0do <= ram0di;
	end else
		ram0do <= ram0[a];
end
always @(posedge sys_clk) begin
	if(we[1]) begin
		ram1[a] <= ram1di;
		ram1do <= ram1di;
	end else
		ram1do <= ram1[a];
end
always @(posedge sys_clk) begin
	if(we[2]) begin
		ram2[a] <= ram2di;
		ram2do <= ram2di;
	end else
		ram2do <= ram2[a];
end
always @(posedge sys_clk) begin
	if(we[3]) begin
		ram3[a] <= ram3di;
		ram3do <= ram3di;
	end else
		ram3do <= ram3[a];
end
always @(posedge sys_clk) begin
	if(we[4]) begin
		ram4[a] <= ram4di;
		ram4do <= ram4di;
	end else
		ram4do <= ram4[a];
end
always @(posedge sys_clk) begin
	if(we[5]) begin
		ram5[a] <= ram5di;
		ram5do <= ram5di;
	end else
		ram5do <= ram5[a];
end
always @(posedge sys_clk) begin
	if(we[6]) begin
		ram6[a] <= ram6di;
		ram6do <= ram6di;
	end else
		ram6do <= ram6[a];
end
always @(posedge sys_clk) begin
	if(we[7]) begin
		ram7[a] <= ram7di;
		ram7do <= ram7di;
	end else
		ram7do <= ram7[a];
end

assign ram0di = di[7:0];
assign ram1di = di[15:8];
assign ram2di = di[23:16];
assign ram3di = di[31:24];
assign ram4di = di[39:32];
assign ram5di = di[47:40];
assign ram6di = di[55:48];
assign ram7di = di[63:56];

assign do = {ram7do, ram6do, ram5do, ram4do, ram3do, ram2do, ram1do, ram0do};

endmodule
